`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   20:50:54 11/08/2018
// Design Name:   Operation5
// Module Name:   /csehome/cobed95/snu-2018-2/LD2018/Assignments/ALU/Operation5Test.v
// Project Name:  ALU
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: Operation5
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module Operation5Test;

	// Inputs
	reg [9:0] operands;

	// Outputs
	wire [6:0] display0;
	wire [6:0] display1;
	wire [6:0] display2;
	wire [6:0] display3;
	wire [6:0] display4;
	wire [6:0] display5;

	// Instantiate the Unit Under Test (UUT)
	Operation5 uut (
		.operands(operands), 
		.display0(display0), 
		.display1(display1), 
		.display2(display2), 
		.display3(display3), 
		.display4(display4), 
		.display5(display5)
	);

	initial begin
		// Initialize Inputs
		operands = 0;

		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here
		operands = 10'b1110100010;
		#100;
		
		operands = 10'b0110100010;
		#100;
		
		operands = 10'b1110100110;
		#100;
		
		operands = 10'b1110100111;
		#100;
		
		operands = 10'b0110100110;
		#100;
		
		operands = 10'b0110100111;
	end
      
endmodule

