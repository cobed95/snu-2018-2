`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   14:43:49 11/07/2018
// Design Name:   Operation1
// Module Name:   /csehome/cobed95/snu-2018-2/LD2018/Assignments/ALU/Operation1Test.v
// Project Name:  ALU
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: Operation1
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module Operation1Test;

	// Inputs
	reg [4:0] operand;

	// Outputs
	wire [6:0] display0;
	wire [6:0] display1;
	wire [6:0] display2;
	wire [6:0] display3;
	wire [6:0] display4;
	wire [6:0] display5;

	// Instantiate the Unit Under Test (UUT)
	Operation1 uut (
		.operand(operand), 
		.display0(display0), 
		.display1(display1), 
		.display2(display2), 
		.display3(display3), 
		.display4(display4), 
		.display5(display5)
	);

	initial begin
		// Initialize Inputs
		operand = 0;

		// Wait 100 ns for global reset to finish
		#20;
      
		// Add stimulus here
		repeat (32) begin 
			operand = operand + 1;
			#20;
		end
		
	end
      
endmodule

